`define VERSION 002