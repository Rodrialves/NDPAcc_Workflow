`define IOB_REVERSE_DATA_W 21
