//Fronte-End
`define IOB_ADDR_W 24
`define IOB_WDATA_W 256
`define IOB_RDATA_W 256
//Back-End
`define BE_ADDR_W 24
`define BE_WDATA_W 256
`define BE_RDATA_W 256