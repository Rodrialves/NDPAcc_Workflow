`define IOB_CACHE_CSRS_ADDR_W 5
`define IOB_CACHE_CSRS_LRU 0
`define IOB_CACHE_CSRS_PLRU_MRU 1
`define IOB_CACHE_CSRS_PLRU_TREE 2
`define IOB_CACHE_CSRS_WRITE_THROUGH 0
`define IOB_CACHE_CSRS_WRITE_BACK 1
`define IOB_CACHE_CSRS_DATA_W 32
`define IOB_CACHE_CSRS_FE_ADDR_W 24
`define IOB_CACHE_CSRS_FE_DATA_W 256
`define IOB_CACHE_CSRS_BE_ADDR_W 24
`define IOB_CACHE_CSRS_BE_DATA_W 256
`define IOB_CACHE_CSRS_NWAYS_W 1
`define IOB_CACHE_CSRS_NLINES_W 10
`define IOB_CACHE_CSRS_WORD_OFFSET_W 3
`define IOB_CACHE_CSRS_WTBUF_DEPTH_W 4
`define IOB_CACHE_CSRS_REP_POLICY 0
`define IOB_CACHE_CSRS_WRITE_POL 0 
`define IOB_CACHE_CSRS_USE_CTRL 0
`define IOB_CACHE_CSRS_USE_CTRL_CNT 0
`define IOB_CACHE_CSRS_VERSION 16'h0002
