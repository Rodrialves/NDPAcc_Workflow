`define IOB_RAM_T2P_HEXFILE "none"
`define IOB_RAM_T2P_ADDR_W 0
`define IOB_RAM_T2P_DATA_W 0
`define IOB_RAM_T2P_MEM_INIT_FILE_INT HEXFILE
