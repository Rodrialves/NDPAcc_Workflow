`define IOB_REG_R_DATA_W 21
`define IOB_REG_R_RST_VAL {DATA_W{1'b0}}
