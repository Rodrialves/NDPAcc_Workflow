`define IOB_REG_DATA_W 1
`define IOB_REG_RST_VAL {DATA_W{1'b0}}
