`timescale 1ns / 1ps
`include "iob_bsp.vh"
`include "iob_cache_aes_ku040_db_g_conf.vh"

module iob_cache_aes_ku040_db_g ();

endmodule
