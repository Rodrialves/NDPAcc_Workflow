`define IOB_REG_RE_DATA_W 21
`define IOB_REG_RE_RST_VAL {DATA_W{1'b0}}
