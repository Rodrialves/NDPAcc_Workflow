`define IOB_REG_E_DATA_W 21
`define IOB_REG_E_RST_VAL {DATA_W{1'b0}}
