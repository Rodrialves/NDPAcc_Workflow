`define IOB_CACHE_SIM_BAUD 3000000
`define IOB_CACHE_SIM_FREQ 100000000
`define IOB_CACHE_SIM_DDR_DATA_W 32
`define IOB_CACHE_SIM_DDR_ADDR_W 24
`define IOB_CACHE_SIM_SIMULATION 1
