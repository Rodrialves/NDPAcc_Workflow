`define IOB_CACHE_AES_KU040_DB_G_BAUD 115200
`define IOB_CACHE_AES_KU040_DB_G_FREQ 100000000
`define IOB_CACHE_AES_KU040_DB_G_DDR_DATA_W 32
`define IOB_CACHE_AES_KU040_DB_G_DDR_ADDR_W 30
`define IOB_CACHE_AES_KU040_DB_G_XILINX 1
