`timescale 1ns / 1ps
`include "iob_bsp.vh"
`include "iob_cache_sim_conf.vh"

module iob_cache_sim ();

endmodule
